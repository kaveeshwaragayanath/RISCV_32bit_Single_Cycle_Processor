module and_gate (
    input logic a,  // Input A
    input logic b,  // Input B
    output logic  y  // Output Y
);

    assign y = a & b;

endmodule
