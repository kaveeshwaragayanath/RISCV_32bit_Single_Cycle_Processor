module ins_memory 
    (input wire clk,          // Clock input
     input wire [7:0] address_in,  
     output wire [31:0] instruction_out  // Data output for read
    );
	 
	  reg [31:0] ins_mem [0:255];
	  
	  assign ins_mem[0]   = 32'b000000000011_01001_010_00110_0000011; //lw             
	  assign ins_mem[4]   = 32'b000000000100_01001_010_00111_0000011; //lw
     assign ins_mem[8]   = 32'b0000000_00111_00110_000_01000_0110011; //add    
     assign ins_mem[12]  = 32'b0100000_00111_00110_000_00011_0110011; //sub  
     assign ins_mem[16]  = 32'b0000000_00111_00110_001_01011_0110011; //sll     
     assign ins_mem[20]  = 32'b0000000_00111_00110_010_01000_0110011; //slt     
     assign ins_mem[24]  = 32'b0000000_00111_00110_011_01111_0110011; //sltu      
     assign ins_mem[28]  = 32'b0000000_00111_00110_100_01011_0110011; // xor     
     assign ins_mem[32]  = 32'b0000000_00111_00110_101_01100_0110011;// srl     
     assign ins_mem[36]  = 32'b0100000_00111_00110_101_01101_0110011;//  sra    
     assign ins_mem[40]  = 32'b0000000_00111_00110_110_01011_0110011;//  or     
     assign ins_mem[44]  = 32'b0000000_00111_00110_111_01111_0110011;// and      
     assign ins_mem[48]  = 32'b0100000_00111_00110_111_01111_0110011;// mul
	  
	  assign ins_mem[52]  = 32'b000000000111_00110_000_00100_0010011;//addi//       
	  assign ins_mem[56]  = 32'b000000010011_00110_010_00100_0010011;//slti
	  assign ins_mem[60]  = 32'b000000010011_00110_011_00100_0010011;//sltiu
	  assign ins_mem[64]  = 32'b000000010011_00110_100_00100_0010011;//xori
	  assign ins_mem[68]  = 32'b000000010011_00110_110_00100_0010011;//ori
	  assign ins_mem[72]  = 32'b000000010011_00110_111_00100_0010011;//andi
	  //
	  assign ins_mem[76]  = 32'b0000010_00111_00110_010_00100_0100011; //sw
	  assign ins_mem[80]  = 32'b0000010_00011_00110_000_00100_0100011; //sb
//	  assign ins_mem[84]  = 32'b0000010_00011_00110_001_00100_0100011; //sh
//	  
//	  //
//	  assign ins_mem[88]  = 32'b000000000011_01001_000_01000_0000011;//lb
//	  assign ins_mem[92]  = 32'b000000000011_01001_001_01000_0000011;//lh
//	  assign ins_mem[96]  = 32'b000000000011_01001_100_01000_0000011;//lbu
//	  assign ins_mem[100]  = 32'b000000000011_01001_101_01000_0000011;//lb
//	  
	  assign ins_mem[84]  = 32'b0000000_01010_00001_000_01000_1100011;//beq
	  assign ins_mem[88]  = 32'b000000000011_01001_000_01000_0000011;//lb
	  assign ins_mem[92]  = 32'b0000000_01001_01010_001_01000_1100011;//bne
	  assign ins_mem[96]  = 32'b000000000011_01001_001_01000_0000011;//lh
	  assign ins_mem[100]  = 32'b0000000_01001_01010_100_01000_1100011;//blt
	  assign ins_mem[104]  = 32'b000000000011_01001_001_01000_0000011;//lh
	  assign ins_mem[108]  = 32'b0000000_01010_01001_101_01000_1100011;//bgt
	  assign ins_mem[112]  = 32'b000000000011_01001_001_01000_0000011;//lh
	  
	  assign ins_mem[116]  = 32'b0000000_01000_00000_000_11000_1101111; //jal
	  assign ins_mem[120]  = 32'b000000000011_01001_001_01000_0000011;//lh
	  assign ins_mem[124]  = 32'b000000000011_01001_001_01000_0000011;//lh
	  
	  
        // Read data from memory at the specified address
     assign    instruction_out = ins_mem[address_in];
    
endmodule 